// Mayu Tatsumi; mtatsumi@g.hmc.edu
// 2025-09-06

module lab2_mt(
	input  logic       reset,
	input  logic [3:0] onboard_s, bboard_s,
	output logic       seg1en, seg2en,
	output logic [4:0] led,
	output logic [6:0] seg
);

// consider adder
// multiplexer
// clk to drive sev-seg outputs (HSOSC required)
// pnp transistors on board for anode

endmodule